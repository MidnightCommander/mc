Tips: Använd C-x t för att kopiera markerade filers namn till kommandoraden.

Tips: Använd C-x p för att kopiera nuvarande katalognamn till kommandoraden.

Tips: Komplettering: anv M-Tab (el Esc+Tab). Tryck två ggr för att få en lista.

Tips: Använd M-p och M-n för att komma åt kommandohistoriken.

Tips: Behöver du skriva ett kontrolltecken? Använd Control-q och tecknet.

Tips: Är du trött på dessa meddelanden? Stäng av dem från Alternativ/Layout-menyn.

Tips: Välja kataloger: Lägg till snedstreck i slutet av det matchande mönstret.

Tips: Om din terminal saknar funktionstangenter, använd ESC+siffersekvens.

Tips: Webbsidan för GNU Midnight Commander: https://midnight-commander.org

Hint: Please file any bug reports at https://github.com/MidnightCommander/mc/issues

Tips: Tab ändrar din nuvarande panel.

Tips: VFS användbarhet: tryck enter på en tar-fil för att se dess innehåll.

Tips: Vi har också en trevlig manualsida.

Tips: Vill du ha navigation i Lynx-stil? Ställ in det i konfigurationsdialogen.

Tips: %-makron fungerar även på kommandoraden.

Tips: M-! tillåter dig att exekvera program och se utskriften i filvisaren.

Tips: Fillistningsformatet kan anpassas; kör "man mc" för detaljer.

Tips: %D/%T expanderar till de markerade filerna i katalogen mitt emot.

Tips: Vill du ha ditt vanliga skal? Tryck C-o och gå tillbaks med C-o igen.

Tips: Att sätta CDPATH-variabeln kan spara tangenttryckningar i cd-kommandon.

Tips: Om du vill se dina .*-filer, ställ in det i konfigurations-dialogen.

Tips: Vill du se dina *~-backupfiler? Ställ in det i konfigurations-dialogen.

Tips: Komplettering funkar på alla inmatningsrutor i dialoger. Tryck på M-Tab.

Tips: På långsamma terminaler kan -s-flaggan hjälpa.

Tips: Sök fil: du kan arbeta med funna filer med panelisera-knappen.

Tips: Vill du göra komplexa sökningar? Använd kommandot Extern panelisering.

Tips: För att ändra katalog under kommandoinmatning, använd M-c (snabb-cd).

Tips: Skalkommandon funkar inte när du är på ett icke-lokalt filsystem.

Tips: Ta tillbaks text från de döda med C-y.

Tips: Fungerar vissa tangenter inte? Se Alternativ/Lär in tangenter.

Tips: för att se utmatningen från ett kommando i filvisaren, använd M-!

Tips: F13 (eller Skift-F3) startar filvisaren i rått läge.

Tips: Du kan specificera editorn för F4 med skalvariabeln EDITOR.

Tips: Du kan välja den externa filvisaren med skalvariabeln VIEWER eller PAGER.

Tips: Du kan slå av alla är-du-säker-frågor i Alternativ/Konfirmation.

Tips: Hoppa till ofta använda kataloger i ett steg med C-\.

Tips: Du kan använda anonym FTP i mc genom att skriva 'cd ftp://dator.se'

Tips: FTP är inbyggt i Midnight Commander, se Fil/FTP-länk-menyn.

Tips: M-t ändrar snabbt listningsläget.

Tips: Du kan specificera användarnamnet med ftps: 'cd ftp://användare@dator.se'

Tips: Du kan bläddra i RPM-filer genom att trycka enter på en RPM-fil.

Tips: För att markera kataloger i markera-dialogrutan, lägg till snedstreck.

Tips: Skift kan behöva hållas ned för att använda klipp och klistra med musen.

Tips: Mata in ofta använda ftp-sajter i favoriter: tryck C-\.
